** Profile: "SCHEMATIC1-TOTO"  [ C:\Users\Sylvain\Desktop\Enseignement_En_Cours\EI\SE3\Ana2\TP\TP2\Ex4\ota-pspicefiles\schematic1\toto.sim ] 

** Creating circuit file "TOTO.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../ota-pspicefiles/ota.lib" 
* From [PSPICE NETLIST] section of C:\Users\Sylvain\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 400u 0 100p 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
